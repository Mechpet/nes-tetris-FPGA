/** font_rom_upscaled:
 * Contains read-only memory pertaining to the text fonts.
 * - Upscaled from an initial 8px by 8px to 16px by 16px.
 * - Tried to preserve the visual style of the font but add smoothness.
 */

module font_rom_upscaled ( input logic [9:0]	addr,
									output logic [15:0]	data
									);

	parameter ADDR_WIDTH = 10;
   parameter DATA_WIDTH =  16;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:735][DATA_WIDTH-1:0] ROM = {
		// Code 0
		16'b0000111111100000, // 0      *******     
		16'b0001111111110000, // 1     *********    
		16'b0011110011111000, // 2    ****  *****   
		16'b0111100001111100, // 3   ****    *****  
		16'b1111000001111110, // 4  ****     ****** 
		16'b1111000011011110, // 5  ****    ** **** 
		16'b1111000110011110, // 6  ****   **  **** 
		16'b1111001100011110, // 7  ****  **   **** 
		16'b1111011000011110, // 8  **** **    **** 
		16'b1111110000011110, // 9  ******     **** 
		16'b1111100000011110, // 10 *****      **** 
		16'b0111110000111100, // 11  *****    ****  
		16'b0011111001111000, // 12   *****  ****   
		16'b0001111111110000, // 13    *********    
		16'b0000111111100000, // 14     *******     
		16'b0000000000000000, // 15                 
		// Code 1
		16'b0000111111100000, // 0      *******     
		16'b0001111111100000, // 1     ********     
		16'b0011111111100000, // 2    *********     
		16'b0011111111100000, // 3    *********     
		16'b0000011111100000, // 4       ******     
		16'b0000011111100000, // 5       ******     
		16'b0000011111100000, // 6       ******     
		16'b0000011111100000, // 7       ******     
		16'b0000011111100000, // 8       ******     
		16'b0000011111100000, // 9       ******     
		16'b0000011111100000, // 10      ******     
		16'b0000011111100000, // 11      ******     
		16'b0000011111100000, // 12      ******     
		16'b0111111111111110, // 13  ************** 
		16'b0111111111111110, // 14  ************** 
		16'b0000000000000000, // 15                 
		// Code 2
		16'b0011111111110000, // 0    **********    
		16'b0111111111111000, // 1   ************   
		16'b1111000000111100, // 2  ****      ****  
		16'b1110000000111100, // 3  ***       ****  
		16'b0000000001111100, // 4           *****  
		16'b0000000011111100, // 5          ******  
		16'b0000000111111100, // 6         *******  
		16'b0000011111111000, // 7       ********   
		16'b0001111111110000, // 8     *********    
		16'b0011111111100000, // 9    *********     
		16'b0111111110000000, // 10  ********       
		16'b1111111000000000, // 11 *******         
		16'b1111110000000000, // 12 ******          
		16'b1111111111111100, // 13 **************  
		16'b1111111111111100, // 14 **************  
		16'b0000000000000000, // 15                 
		// Code 3
		16'b0011111111111110, // 0    ************* 
		16'b0011111111111110, // 1    ************* 
		16'b0000000001111100, // 2           *****  
		16'b0000000011111000, // 3          *****   
		16'b0000000111110000, // 4         *****    
		16'b0000001111100000, // 5        *****     
		16'b0000011111111000, // 6       ********   
		16'b0000111111111100, // 7      **********  
		16'b0000111111111110, // 8      *********** 
		16'b0000000000111110, // 9            ***** 
		16'b0000000000011110, // 10            **** 
		16'b1111000000011110, // 11 ****       **** 
		16'b1111100000111110, // 12 *****     ***** 
		16'b0111111111111100, // 13  *************  
		16'b0011111111111000, // 14   ***********   
		16'b0000000000000000, // 15                 
		// Code 4
		16'b0000001111111000, // 0        *******   
		16'b0000011111111000, // 1       ********   
		16'b0000111111111000, // 2      *********   
		16'b0001111111111000, // 3     **********   
		16'b0011111001111000, // 4    *****  ****   
		16'b0111110001111000, // 5   *****   ****   
		16'b1111100001111000, // 6  *****    ****   
		16'b1111000001111000, // 7  ****     ****   
		16'b1111000001111000, // 8  ****     ****   
		16'b1111111111111110, // 9  *************** 
		16'b1111111111111110, // 10 *************** 
		16'b0000000001111000, // 11          ****   
		16'b0000000001111000, // 12          ****   
		16'b0000000001111000, // 13          ****   
		16'b0000000001111000, // 14          ****   
		16'b0000000000000000, // 15                 
		// Code 5
		16'b1111111111111100, // 0  **************  
		16'b1111111111111100, // 1  **************  
		16'b1111100000000000, // 2  *****           
		16'b1111100000000000, // 3  *****           
		16'b1111111111100000, // 4  ***********     
		16'b1111111111110000, // 5  ************    
		16'b1111111111111000, // 6  *************   
		16'b0000000111111100, // 7         *******  
		16'b0000000011111100, // 8          ******  
		16'b0000000001111100, // 9           *****  
		16'b0000000001111100, // 10          *****  
		16'b1111000001111100, // 11 ****     *****  
		16'b1111100011111100, // 12 *****   ******  
		16'b0111111111111000, // 13  ************   
		16'b0011111111100000, // 14   *********     
		16'b0000000000000000, // 15                 
		// Code 6
		16'b0000111111111000, // 0      *********   
		16'b0001111111111000, // 1     **********   
		16'b0011111000000000, // 2    *****         
		16'b0111110000000000, // 3   *****          
		16'b1111100000000000, // 4  *****           
		16'b1111000000000000, // 5  ****            
		16'b1111111111111000, // 6  *************   
		16'b1111111111111100, // 7  **************  
		16'b1111111111111100, // 8  **************  
		16'b1111100000111110, // 9  *****     ***** 
		16'b1111000000011110, // 10 ****       **** 
		16'b1111000000011110, // 11 ****       **** 
		16'b1111100000111110, // 12 *****     ***** 
		16'b0111111111111100, // 13  *************  
		16'b0011111111111000, // 14   ***********   
		16'b0000000000000000, // 15                 
		// Code 7
		16'b0111111111111110, // 0   ************** 
		16'b1111111111111110, // 1  *************** 
		16'b1111000000011110, // 2  ****       **** 
		16'b1111000000111110, // 3  ****      ***** 
		16'b0000000001111100, // 4           *****  
		16'b0000000011111000, // 5          *****   
		16'b0000000111110000, // 6         *****    
		16'b0000001111100000, // 7        *****     
		16'b0000011111100000, // 8       ******     
		16'b0000011111000000, // 9       *****      
		16'b0000111111000000, // 10     ******      
		16'b0000111110000000, // 11     *****       
		16'b0000111110000000, // 12     *****       
		16'b0000111110000000, // 13     *****       
		16'b0000111110000000, // 14     *****       
		16'b0000000000000000, // 15                 
		// Code 8
		16'b0011111111100000, // 0    *********     
		16'b0111111111110000, // 1   ***********    
		16'b1111000000111000, // 2  ****      ***   
		16'b1111000000011000, // 3  ****       **   
		16'b1111100000011000, // 4  *****      **   
		16'b0111110000011000, // 5   *****     **   
		16'b0011111111110000, // 6    **********    
		16'b0011111111100000, // 7    *********     
		16'b0111111111111000, // 8   ************   
		16'b1110001111111100, // 9  ***   ********  
		16'b1100000011111110, // 10 **      ******* 
		16'b1100000000111110, // 11 **        ***** 
		16'b1110000000011110, // 12 ***        **** 
		16'b0111111111111100, // 13  *************  
		16'b0011111111111000, // 14   ***********   
		16'b0000000000000000, // 15                 
		// Code 9
		16'b0011111111111000, // 0    ***********   
		16'b0111111111111100, // 1   *************  
		16'b1111100000111110, // 2  *****     ***** 
		16'b1111000000011110, // 3  ****       **** 
		16'b1111000000011110, // 4  ****       **** 
		16'b1111100000111110, // 5  *****     ***** 
		16'b0111111111111110, // 6   ************** 
		16'b0111111111111110, // 7   ************** 
		16'b0011111111111110, // 8    ************* 
		16'b0000000000011110, // 9             **** 
		16'b0000000000111110, // 10           ***** 
		16'b0000000001111100, // 11          *****  
		16'b0000000011111000, // 12         *****   
		16'b0011111111110000, // 13   **********    
		16'b0011111111100000, // 14   *********     
		16'b0000000000000000, // 15                 
		// Code 10
		16'b0000111111100000, // 0      *******     
		16'b0001111111110000, // 1     *********    
		16'b0011111111111000, // 2    ***********   
		16'b0111110001111100, // 3   *****   *****  
		16'b1111100000111110, // 4  *****     ***** 
		16'b1111000000011110, // 5  ****       **** 
		16'b1111000000011110, // 6  ****       **** 
		16'b1111000000011110, // 7  ****       **** 
		16'b1111000000011110, // 8  ****       **** 
		16'b1111111111111110, // 9  *************** 
		16'b1111111111111110, // 10 *************** 
		16'b1111000000011110, // 11 ****       **** 
		16'b1111000000011110, // 12 ****       **** 
		16'b1111000000011110, // 13 ****       **** 
		16'b1111000000011110, // 14 ****       **** 
		16'b0000000000000000, // 15                 
		// Code 11
		16'b1111111111111000, // 0  *************   
		16'b1111111111111100, // 1  **************  
		16'b1111000000111110, // 2  ****      ***** 
		16'b1111000000011110, // 3  ****       **** 
		16'b1111000000011110, // 4  ****       **** 
		16'b1111000000111110, // 5  ****      ***** 
		16'b1111111111111100, // 6  **************  
		16'b1111111111111000, // 7  *************   
		16'b1111111111111100, // 8  **************  
		16'b1111000000111110, // 9  ****      ***** 
		16'b1111000000011110, // 10 ****       **** 
		16'b1111000000011110, // 11 ****       **** 
		16'b1111000000111110, // 12 ****      ***** 
		16'b1111111111111100, // 13 **************  
		16'b1111111111111000, // 14 *************   
		16'b0000000000000000, // 15                 
		// Code 12
		16'b0000111111111000, // 0      *********   
		16'b0001111111111100, // 1     ***********  
		16'b0011111000111110, // 2    *****   ***** 
		16'b0111110000011110, // 3   *****     **** 
		16'b1111100000000000, // 4  *****           
		16'b1111000000000000, // 5  ****            
		16'b1111000000000000, // 6  ****            
		16'b1111000000000000, // 7  ****            
		16'b1111000000000000, // 8  ****            
		16'b1111000000000000, // 9  ****            
		16'b1111100000000000, // 10 *****           
		16'b0111110000011110, // 11  *****     **** 
		16'b0011111000111110, // 12   *****   ***** 
		16'b0001111111111100, // 13    ***********  
		16'b0000111111111000, // 14     *********   
		16'b0000000000000000, // 15                 
		// Code 13
		16'b1111111111100000, // 0  ***********     
		16'b1111111111110000, // 1  ************    
		16'b1111000011111000, // 2  ****    *****   
		16'b1111000001111100, // 3  ****     *****  
		16'b1111000000111110, // 4  ****      ***** 
		16'b1111000000011110, // 5  ****       **** 
		16'b1111000000011110, // 6  ****       **** 
		16'b1111000000011110, // 7  ****       **** 
		16'b1111000000011110, // 8  ****       **** 
		16'b1111000000011110, // 9  ****       **** 
		16'b1111000000111110, // 10 ****      ***** 
		16'b1111000001111100, // 11 ****     *****  
		16'b1111000011111000, // 12 ****    *****   
		16'b1111111111110000, // 13 ************    
		16'b1111111111100000, // 14 ***********     
		16'b0000000000000000, // 15                 
		// Code 14
		16'b1111111111111110, // 0  *************** 
		16'b1111111111111110, // 1  *************** 
		16'b1111000000000000, // 2  ****            
		16'b1111000000000000, // 3  ****            
		16'b1111000000000000, // 4  ****            
		16'b1111000000000000, // 5  ****            
		16'b1111111111111000, // 6  *************   
		16'b1111111111111000, // 7  *************   
		16'b1111111111111000, // 8  *************   
		16'b1111000000000000, // 9  ****            
		16'b1111000000000000, // 10 ****            
		16'b1111000000000000, // 11 ****            
		16'b1111000000000000, // 12 ****            
		16'b1111111111111110, // 13 *************** 
		16'b1111111111111110, // 14 *************** 
		16'b0000000000000000, // 15                 
		// Code 15
		16'b1111111111111110, // 0  *************** 
		16'b1111111111111110, // 1  *************** 
		16'b1111000000000000, // 2  ****            
		16'b1111000000000000, // 3  ****            
		16'b1111000000000000, // 4  ****            
		16'b1111000000000000, // 5  ****            
		16'b1111111111111000, // 6  *************   
		16'b1111111111111000, // 7  *************   
		16'b1111111111111000, // 8  *************   
		16'b1111000000000000, // 9  ****            
		16'b1111000000000000, // 10 ****            
		16'b1111000000000000, // 11 ****            
		16'b1111000000000000, // 12 ****            
		16'b1111000000000000, // 13 ****            
		16'b1111000000000000, // 14 ****            
		16'b0000000000000000, // 15                 
		// Code 16
		16'b0000111111111110, // 0      *********** 
		16'b0001111111111110, // 1     ************ 
		16'b0011111000000000, // 2    *****         
		16'b0111110000000000, // 3   *****          
		16'b1111100000000000, // 4  *****           
		16'b1111000000000000, // 5  ****            
		16'b1111000001111110, // 6  ****     ****** 
		16'b1111000001111110, // 7  ****     ****** 
		16'b1111000001111110, // 8  ****     ****** 
		16'b1111000000011110, // 9  ****       **** 
		16'b1111100000011110, // 10 *****      **** 
		16'b0111110000011110, // 11  *****     **** 
		16'b0011111000011110, // 12   *****    **** 
		16'b0001111111111110, // 13    ************ 
		16'b0000111111111110, // 14     *********** 
		16'b0000000000000000, // 15                 
		// Code 17
		16'b1111000000011110, // 0  ****       **** 
		16'b1111000000011110, // 1  ****       **** 
		16'b1111000000011110, // 2  ****       **** 
		16'b1111000000011110, // 3  ****       **** 
		16'b1111000000011110, // 4  ****       **** 
		16'b1111000000011110, // 5  ****       **** 
		16'b1111111111111110, // 6  *************** 
		16'b1111111111111110, // 7  *************** 
		16'b1111111111111110, // 8  *************** 
		16'b1111000000011110, // 9  ****       **** 
		16'b1111000000011110, // 10 ****       **** 
		16'b1111000000011110, // 11 ****       **** 
		16'b1111000000011110, // 12 ****       **** 
		16'b1111000000011110, // 13 ****       **** 
		16'b1111000000011110, // 14 ****       **** 
		16'b0000000000000000, // 15                 
		// Code 18
		16'b0111111111111110, // 0   ************** 
		16'b0111111111111110, // 1   ************** 
		16'b0000011111100000, // 2       ******     
		16'b0000011111100000, // 3       ******     
		16'b0000011111100000, // 4       ******     
		16'b0000011111100000, // 5       ******     
		16'b0000011111100000, // 6       ******     
		16'b0000011111100000, // 7       ******     
		16'b0000011111100000, // 8       ******     
		16'b0000011111100000, // 9       ******     
		16'b0000011111100000, // 10      ******     
		16'b0000011111100000, // 11      ******     
		16'b0000011111100000, // 12      ******     
		16'b0111111111111110, // 13  ************** 
		16'b0111111111111110, // 14  ************** 
		16'b0000000000000000, // 15                 
		// Code 19
		16'b0000000000011110, // 0             **** 
		16'b0000000000011110, // 1             **** 
		16'b0000000000011110, // 2             **** 
		16'b0000000000011110, // 3             **** 
		16'b0000000000011110, // 4             **** 
		16'b0000000000011110, // 5             **** 
		16'b0000000000011110, // 6             **** 
		16'b0000000000011110, // 7             **** 
		16'b0000000000011110, // 8             **** 
		16'b0000000000011110, // 9             **** 
		16'b0000000000011110, // 10            **** 
		16'b1111000000011110, // 11 ****       **** 
		16'b1111100000111110, // 12 *****     ***** 
		16'b0111111111111100, // 13  *************  
		16'b0011111111111000, // 14   ***********   
		16'b0000000000000000, // 15                 
		// Code 20
		16'b1111100000111110, // 0  *****     ***** 
		16'b1111100001111110, // 1  *****    ****** 
		16'b1111100011111100, // 2  *****   ******  
		16'b1111100111111000, // 3  *****  ******   
		16'b1111101111110000, // 4  ***** ******    
		16'b1111111111100000, // 5  ***********     
		16'b1111111111000000, // 6  **********      
		16'b1111111110000000, // 7  *********       
		16'b1111111110000000, // 8  *********       
		16'b1111111111000000, // 9  **********      
		16'b1111111111100000, // 10 ***********     
		16'b1111111111110000, // 11 ************    
		16'b1111100111111000, // 12 *****  ******   
		16'b1111100011111100, // 13 *****   ******  
		16'b1111100001111110, // 14 *****    ****** 
		16'b0000000000000000, // 15                 
		// Code 21
		16'b1111000000000000, // 0  ****            
		16'b1111000000000000, // 1  ****            
		16'b1111000000000000, // 2  ****            
		16'b1111000000000000, // 3  ****            
		16'b1111000000000000, // 4  ****            
		16'b1111000000000000, // 5  ****            
		16'b1111000000000000, // 6  ****            
		16'b1111000000000000, // 7  ****            
		16'b1111000000000000, // 8  ****            
		16'b1111000000000000, // 9  ****            
		16'b1111000000000000, // 10 ****            
		16'b1111000000000000, // 11 ****            
		16'b1111111111111110, // 12 *************** 
		16'b1111111111111110, // 13 *************** 
		16'b1111111111111110, // 14 *************** 
		16'b0000000000000000, // 15                 
		// Code 22
		16'b1111000000011110, // 0  ****       **** 
		16'b1111100000111110, // 1  *****     ***** 
		16'b1111110001111110, // 2  ******   ****** 
		16'b1111111011111110, // 3  ******* ******* 
		16'b1111111111111110, // 4  *************** 
		16'b1111111111111110, // 5  *************** 
		16'b1111111111111110, // 6  *************** 
		16'b1111111111111110, // 7  *************** 
		16'b1111111111111110, // 8  *************** 
		16'b1111011111011110, // 9  **** ***** **** 
		16'b1111001110011110, // 10 ****  ***  **** 
		16'b1111000100011110, // 11 ****   *   **** 
		16'b1111000000011110, // 12 ****       **** 
		16'b1111000000011110, // 13 ****       **** 
		16'b1111000000011110, // 14 ****       **** 
		16'b0000000000000000, // 15                 
		// Code 23
		16'b1111100000011110, // 0  *****      **** 
		16'b1111110000011110, // 1  ******     **** 
		16'b1111111000011110, // 2  *******    **** 
		16'b1111111100011110, // 3  ********   **** 
		16'b1111111110011110, // 4  *********  **** 
		16'b1111111111011110, // 5  ********** **** 
		16'b1111111111111110, // 6  *************** 
		16'b1111111111111110, // 7  *************** 
		16'b1111111111111110, // 8  *************** 
		16'b1111011111111110, // 9  **** ********** 
		16'b1111001111111110, // 10 ****  ********* 
		16'b1111000111111110, // 11 ****   ******** 
		16'b1111000011111110, // 12 ****    ******* 
		16'b1111000001111110, // 13 ****     ****** 
		16'b1111000000111110, // 14 ****      ***** 
		16'b0000000000000000, // 15                 
		// Code 24
		16'b0011111111111000, // 0    ***********   
		16'b0111111111111100, // 1   *************  
		16'b1111100000111110, // 2  *****     ***** 
		16'b1111000000011110, // 3  ****       **** 
		16'b1111000000011110, // 4  ****       **** 
		16'b1111000000011110, // 5  ****       **** 
		16'b1111000000011110, // 6  ****       **** 
		16'b1111000000011110, // 7  ****       **** 
		16'b1111000000011110, // 8  ****       **** 
		16'b1111000000011110, // 9  ****       **** 
		16'b1111000000011110, // 10 ****       **** 
		16'b1111000000011110, // 11 ****       **** 
		16'b1111100000111110, // 12 *****     ***** 
		16'b0111111111111100, // 13  *************  
		16'b0011111111111000, // 14   ***********   
		16'b0000000000000000, // 15                 
		// Code 25
		16'b1111111111111000, // 0  *************   
		16'b1111111111111100, // 1  **************  
		16'b1111000000111110, // 2  ****      ***** 
		16'b1111000000011110, // 3  ****       **** 
		16'b1111000000011110, // 4  ****       **** 
		16'b1111000000011110, // 5  ****       **** 
		16'b1111000000011110, // 6  ****       **** 
		16'b1111000000011110, // 7  ****       **** 
		16'b1111000000111110, // 8  ****      ***** 
		16'b1111111111111100, // 9  **************  
		16'b1111111111111000, // 10 *************   
		16'b1111000000000000, // 11 ****            
		16'b1111000000000000, // 12 ****            
		16'b1111000000000000, // 13 ****            
		16'b1111000000000000, // 14 ****            
		16'b0000000000000000, // 15                 
		// Code 26
		16'b0011111111111000, // 0    ***********   
		16'b0111111111111100, // 1   *************  
		16'b1111100000111110, // 2  *****     ***** 
		16'b1111000000011110, // 3  ****       **** 
		16'b1111000000011110, // 4  ****       **** 
		16'b1111000000011110, // 5  ****       **** 
		16'b1111000000011110, // 6  ****       **** 
		16'b1111000000011110, // 7  ****       **** 
		16'b1111000111111110, // 8  ****   ******** 
		16'b1111000111111110, // 9  ****   ******** 
		16'b1111000011111100, // 10 ****    ******  
		16'b1111000001111000, // 11 ****     ****   
		16'b1111100011111100, // 12 *****   ******  
		16'b0111111111101110, // 13  ********** *** 
		16'b0011111111000110, // 14   ********   ** 
		16'b0000000000000000, // 15                 
		// Code 27
		16'b1111111111110000, // 0  ************    
		16'b1111111111111000, // 1  *************   
		16'b1111000001111100, // 2  ****     *****  
		16'b1111000000111110, // 3  ****      ***** 
		16'b1111000000011110, // 4  ****       **** 
		16'b1111000000011110, // 5  ****       **** 
		16'b1111000000111110, // 6  ****      ***** 
		16'b1111000001111100, // 7  ****     *****  
		16'b1111111111111000, // 8  *************   
		16'b1111111111110000, // 9  ************    
		16'b1111111111100000, // 10 ***********     
		16'b1111001111110000, // 11 ****  ******    
		16'b1111000111111000, // 12 ****   ******   
		16'b1111000011111100, // 13 ****    ******  
		16'b1111000001111110, // 14 ****     ****** 
		16'b0000000000000000, // 15                 
		// Code 28
		16'b0011111111100000, // 0    *********     
		16'b0111111111110000, // 1   ***********    
		16'b1111100011111000, // 2  *****   *****   
		16'b1111000001111000, // 3  ****     ****   
		16'b1111000000000000, // 4  ****            
		16'b1111100000000000, // 5  *****           
		16'b0111111111110000, // 6   ***********    
		16'b0011111111111000, // 7    ***********   
		16'b0001111111111100, // 8     ***********  
		16'b0000000000111110, // 9            ***** 
		16'b0000000000011110, // 10            **** 
		16'b1111000000011110, // 11 ****       **** 
		16'b1111100000111110, // 12 *****     ***** 
		16'b0111111111111100, // 13  *************  
		16'b0011111111111000, // 14   ***********   
		16'b0000000000000000, // 15                 
		// Code 29
		16'b0111111111111110, // 0   ************** 
		16'b0111111111111110, // 1   ************** 
		16'b0000011111100000, // 2       ******     
		16'b0000011111100000, // 3       ******     
		16'b0000011111100000, // 4       ******     
		16'b0000011111100000, // 5       ******     
		16'b0000011111100000, // 6       ******     
		16'b0000011111100000, // 7       ******     
		16'b0000011111100000, // 8       ******     
		16'b0000011111100000, // 9       ******     
		16'b0000011111100000, // 10      ******     
		16'b0000011111100000, // 11      ******     
		16'b0000011111100000, // 12      ******     
		16'b0000011111100000, // 13      ******     
		16'b0000011111100000, // 14      ******     
		16'b0000000000000000, // 15                 
		// Code 30
		16'b1111000000011110, // 0  ****       **** 
		16'b1111000000011110, // 1  ****       **** 
		16'b1111000000011110, // 2  ****       **** 
		16'b1111000000011110, // 3  ****       **** 
		16'b1111000000011110, // 4  ****       **** 
		16'b1111000000011110, // 5  ****       **** 
		16'b1111000000011110, // 6  ****       **** 
		16'b1111000000011110, // 7  ****       **** 
		16'b1111000000011110, // 8  ****       **** 
		16'b1111000000011110, // 9  ****       **** 
		16'b1111000000011110, // 10 ****       **** 
		16'b1111000000011110, // 11 ****       **** 
		16'b1111100000111110, // 12 *****     ***** 
		16'b0111111111111100, // 13  *************  
		16'b0011111111111000, // 14   ***********   
		16'b0000000000000000, // 15                 
		// Code 31
		16'b1111000000011110, // 0  ****       **** 
		16'b1111000000011110, // 1  ****       **** 
		16'b1111000000011110, // 2  ****       **** 
		16'b1111000000011110, // 3  ****       **** 
		16'b1111000000011110, // 4  ****       **** 
		16'b1111100000111110, // 5  *****     ***** 
		16'b1111100000111110, // 6  *****     ***** 
		16'b1111110001111110, // 7  ******   ****** 
		16'b1111111011111110, // 8  ******* ******* 
		16'b0111111111111100, // 9   *************  
		16'b0011111111111000, // 10   ***********   
		16'b0001111111110000, // 11    *********    
		16'b0000111111100000, // 12     *******     
		16'b0000011111000000, // 13      *****      
		16'b0000001110000000, // 14       ***       
		16'b0000000000000000, // 15                 
		// Code 32
		16'b1111000000011110, // 0  ****       **** 
		16'b1111000000011110, // 1  ****       **** 
		16'b1111000000011110, // 2  ****       **** 
		16'b1111000100011110, // 3  ****   *   **** 
		16'b1111001110011110, // 4  ****  ***  **** 
		16'b1111011111011110, // 5  **** ***** **** 
		16'b1111111111111110, // 6  *************** 
		16'b1111111111111110, // 7  *************** 
		16'b1111111111111110, // 8  *************** 
		16'b1111111111111110, // 9  *************** 
		16'b1111111111111110, // 10 *************** 
		16'b1111111011111110, // 11 ******* ******* 
		16'b1111110001111110, // 12 ******   ****** 
		16'b1111100000111110, // 13 *****     ***** 
		16'b1111000000011110, // 14 ****       **** 
		16'b0000000000000000, // 15                 
		// Code 33
		16'b1111000000011110, // 0  ****       **** 
		16'b1111100000111110, // 1  *****     ***** 
		16'b1111110001111110, // 2  ******   ****** 
		16'b1111111011111110, // 3  ******* ******* 
		16'b0111111111111100, // 4   *************  
		16'b0011111111111000, // 5    ***********   
		16'b0001111111110000, // 6     *********    
		16'b0000111111100000, // 7      *******     
		16'b0001111111110000, // 8     *********    
		16'b0011111111111000, // 9    ***********   
		16'b0111111111111100, // 10  *************  
		16'b1111111011111110, // 11 ******* ******* 
		16'b1111110001111110, // 12 ******   ****** 
		16'b1111100000111110, // 13 *****     ***** 
		16'b1111000000011110, // 14 ****       **** 
		16'b0000000000000000, // 15                 
		// Code 34
		16'b0111100000011110, // 0   ****      **** 
		16'b0111100000011110, // 1   ****      **** 
		16'b0111100000011110, // 2   ****      **** 
		16'b0111100000011110, // 3   ****      **** 
		16'b0111100000011110, // 4   ****      **** 
		16'b0111110000111110, // 5   *****    ***** 
		16'b0011111111111100, // 6    ************  
		16'b0001111111111000, // 7     **********   
		16'b0001111111111000, // 8     **********   
		16'b0000111111110000, // 9      ********    
		16'b0000011111100000, // 10      ******     
		16'b0000011111100000, // 11      ******     
		16'b0000011111100000, // 12      ******     
		16'b0000011111100000, // 13      ******     
		16'b0000011111100000, // 14      ******     
		16'b0000000000000000, // 15                 
		// Code 35
		16'b1111111111111110, // 0  *************** 
		16'b1111111111111110, // 1  *************** 
		16'b0000000001111110, // 2           ****** 
		16'b0000000011111110, // 3          ******* 
		16'b0000000111111100, // 4         *******  
		16'b0000001111111000, // 5        *******   
		16'b0000011111110000, // 6       *******    
		16'b0000111111100000, // 7      *******     
		16'b0001111111000000, // 8     *******      
		16'b0011111110000000, // 9    *******       
		16'b0111111100000000, // 10  *******        
		16'b1111111000000000, // 11 *******         
		16'b1111110000000000, // 12 ******          
		16'b1111111111111110, // 13 *************** 
		16'b1111111111111110, // 14 *************** 
		16'b0000000000000000, // 15                 
		// Code 36
		16'b0000000000000000, // 0                  
		16'b0000000000000000, // 1                  
		16'b0000000000000000, // 2                  
		16'b0000000000000000, // 3                  
		16'b0000000000000000, // 4                  
		16'b0000000000000000, // 5                  
		16'b0000000000000000, // 6                  
		16'b0000000000000000, // 7                  
		16'b0000000000000000, // 8                  
		16'b0000000000000000, // 9                  
		16'b0000000000000000, // 10                 
		16'b0011110000000000, // 11   ****          
		16'b0011110000000000, // 12   ****          
		16'b0011110000000000, // 13   ****          
		16'b0011110000000000, // 14   ****          
		16'b0000000000000000, // 15                 
		// Code 37
		16'b0000000000000000, // 0                  
		16'b0000000000000000, // 1                  
		16'b0000000000000000, // 2                  
		16'b0000000000000000, // 3                  
		16'b0000000000000000, // 4                  
		16'b0000000000000000, // 5                  
		16'b0000000000000000, // 6                  
		16'b0000000000000000, // 7                  
		16'b0000000000000000, // 8                  
		16'b0000000000000000, // 9                  
		16'b0000001111000000, // 10       ****      
		16'b0000001111000000, // 11       ****      
		16'b0000000011000000, // 12         **      
		16'b0000000011000000, // 13         **      
		16'b0000001100000000, // 14       **        
		16'b0000001100000000, // 15       **        
		// Code 38
		16'b0000011111100000, // 0       ******     
		16'b0000011111100000, // 1       ******     
		16'b0000011111100000, // 2       ******     
		16'b0000011111100000, // 3       ******     
		16'b0000011111100000, // 4       ******     
		16'b0000011111100000, // 5       ******     
		16'b0000011111100000, // 6       ******     
		16'b0000011111100000, // 7       ******     
		16'b0000011111100000, // 8       ******     
		16'b0000011111100000, // 9       ******     
		16'b0000011111100000, // 10      ******     
		16'b0000000000000000, // 11                 
		16'b0000000000000000, // 12                 
		16'b0000011111100000, // 13      ******     
		16'b0000011111100000, // 14      ******     
		16'b0000000000000000, // 15                 
		// Code 39
		16'b0000110000110000, // 0      **    **    
		16'b0000110000110000, // 1      **    **    
		16'b0011111111111100, // 2    ************  
		16'b0011111111111100, // 3    ************  
		16'b0000110000110000, // 4      **    **    
		16'b0000110000110000, // 5      **    **    
		16'b0000110000110000, // 6      **    **    
		16'b0000110000110000, // 7      **    **    
		16'b0000110000110000, // 8      **    **    
		16'b0011111111111100, // 9    ************  
		16'b0011111111111100, // 10   ************  
		16'b0000110000110000, // 11     **    **    
		16'b0000110000110000, // 12     **    **    
		16'b0000000000000000, // 13                 
		16'b0000000000000000, // 14                 
		16'b0000000000000000, // 15                 
		// Code 40
		16'b0000000000000000, // 0                  
		16'b0000000000000000, // 1                  
		16'b0000000000000000, // 2                  
		16'b0000000000000000, // 3                  
		16'b0000000000000000, // 4                  
		16'b0000000000000000, // 5                  
		16'b0000000000000000, // 6                  
		16'b0011111111111100, // 7    ************  
		16'b0011111111111100, // 8    ************  
		16'b0011111111111100, // 9    ************  
		16'b0000000000000000, // 10                 
		16'b0000000000000000, // 11                 
		16'b0000000000000000, // 12                 
		16'b0000000000000000, // 13                 
		16'b0000000000000000, // 14                 
		16'b0000000000000000, // 15                 
		// Code 41
		16'b0000000000001111, // 0              ****
		16'b0000000000011111, // 1             *****
		16'b0000000000111110, // 2            ***** 
		16'b0000000001111100, // 3           *****  
		16'b0000000011111000, // 4          *****   
		16'b0000000111110000, // 5         *****    
		16'b0000001111100000, // 6        *****     
		16'b0000011111000000, // 7       *****      
		16'b0000111110000000, // 8      *****       
		16'b0001111100000000, // 9     *****        
		16'b0011111000000000, // 10   *****         
		16'b0111110000000000, // 11  *****          
		16'b1111100000000000, // 12 *****           
		16'b1111000000000000, // 13 ****            
		16'b0000000000000000, // 14                 
		16'b0000000000000000, // 15                 
		// Code 42
		16'b0000000000000000, // 0                  
		16'b0000000000000000, // 1                  
		16'b0000001111000000, // 2        ****      
		16'b0000001111000000, // 3        ****      
		16'b0000001111000000, // 4        ****      
		16'b0000001111000000, // 5        ****      
		16'b0000000000000000, // 6                  
		16'b0000000000000000, // 7                  
		16'b0000000000000000, // 8                  
		16'b0000000000000000, // 9                  
		16'b0000001111000000, // 10       ****      
		16'b0000001111000000, // 11       ****      
		16'b0000001111000000, // 12       ****      
		16'b0000001111000000, // 13       ****      
		16'b0000000000000000, // 14                 
		16'b0000000000000000, // 15                 
		// Code 43
		16'b0000000000000000, // 0                  
		16'b0000000000000000, // 1                  
		16'b0000000000000000, // 2                  
		16'b0000000000000000, // 3                  
		16'b0011111111111100, // 4    ************  
		16'b0011111111111100, // 5    ************  
		16'b0000000000000000, // 6                  
		16'b0000000000000000, // 7                  
		16'b0000000000000000, // 8                  
		16'b0000000000000000, // 9                  
		16'b0011111111111100, // 10   ************  
		16'b0011111111111100, // 11   ************  
		16'b0000000000000000, // 12                 
		16'b0000000000000000, // 13                 
		16'b0000000000000000, // 14                 
		16'b0000000000000000, // 15                 
		// Code 44
		16'b0000111111110000, // 0      ********    
		16'b0001111111111000, // 1     **********   
		16'b0011100000011100, // 2    ***      ***  
		16'b0111000000001110, // 3   ***        *** 
		16'b1110001111000111, // 4  ***   ****   ***
		16'b1100011111100011, // 5  **   ******   **
		16'b1100011001100011, // 6  **   **  **   **
		16'b1100011000000011, // 7  **   **       **
		16'b1100011000000011, // 8  **   **       **
		16'b1100011001100011, // 9  **   **  **   **
		16'b1100011111100011, // 10 **   ******   **
		16'b1110001111000111, // 11 ***   ****   ***
		16'b0111000000001110, // 12  ***        *** 
		16'b0011100000011100, // 13   ***      ***  
		16'b0001111111111000, // 14    **********   
		16'b0000111111110000, // 15     ********    
		// Code 45
		16'b0000000000000000, // 0                  
		16'b0000000000000000, // 1                  
		16'b0000000000000000, // 2                  
		16'b0000000000000000, // 3                  
		16'b0000000000000000, // 4                  
		16'b0000000000000000, // 5                  
		16'b0000000000000000, // 6                  
		16'b0000000000000000, // 7                  
		16'b0000000000000000, // 8                  
		16'b0000000000000000, // 9                  
		16'b0000000000000000, // 10                 
		16'b0000000000000000, // 11                 
		16'b0000000000000000, // 12                 
		16'b0000000000000000, // 13                 
		16'b0000000000000000, // 14                 
		16'b0000000000000000  // 15                         
	};
	assign data = ROM[addr];
endmodule  