package my_pkg;

parameter [6:0] score_label_left_col = 68;
parameter [6:0] score_label_right_col = 72;
parameter [6:0] score_label_row = 12;
parameter [9:0] start_S = 6'h1C * 8;
parameter [9:0] start_C = 6'h0C * 8;
parameter [9:0] start_O = 6'h18 * 8;
parameter [9:0] start_R = 6'h1B * 8;
parameter [9:0] start_E = 6'h0E * 8;

endpackage