module font_rom ( input [5:0]	addr,
						output [7:0]	data
					 );

	parameter ADDR_WIDTH = 6;
   parameter DATA_WIDTH =  8;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
			// code x00
        8'b00111000, // 0   ***   
        8'b01001100, // 1  *  **  
        8'b11000110, // 2 **   ** 
        8'b11000110, // 3 **   ** 
        8'b11000110, // 4 **   ** 
        8'b01100100, // 5  **  *  
        8'b00111000, // 6   ***   
        8'b00000000, // 7         
         // code x01
        8'b00110000, // 0   **    
        8'b01110000, // 1  ***    
        8'b00110000, // 2   **    
        8'b00110000, // 3   **    
        8'b00110000, // 4   **    
        8'b00110000, // 5   **    
        8'b11111100, // 6 ******  
        8'b00000000, // 7         
         // code x02
        8'b01111100, // 0  *****  
        8'b11000110, // 1 **   ** 
        8'b00001110, // 2     *** 
        8'b00011110, // 3    **** 
        8'b00111100, // 4   ****  
        8'b11100000, // 5 ***     
        8'b11111110, // 6 ******* 
        8'b00000000, // 7         
         // code x03
        8'b01111110, // 0  ****** 
        8'b00001100, // 1     **  
        8'b00011000, // 2    **   
        8'b00111100, // 3   ****  
        8'b00000110, // 4      ** 
        8'b11000110, // 5 **   ** 
        8'b01111100, // 6  *****  
        8'b00000000, // 7         
         // code x04
        8'b00011100, // 0    ***  
        8'b00111100, // 1   ****  
        8'b01101100, // 2  ** **  
        8'b11001100, // 3 **  **  
        8'b11111110, // 4 ******* 
        8'b00001100, // 5     **  
        8'b00001100, // 6     **  
        8'b00000000, // 7         
         // code x05
        8'b11111100, // 0 ******  
        8'b11000000, // 1 **      
        8'b11111100, // 2 ******  
        8'b00000110, // 3      ** 
        8'b00000110, // 4      ** 
        8'b11000110, // 5 **   ** 
        8'b01111100, // 6  *****  
        8'b00000000, // 7         
         // code x06
        8'b00111100, // 0   ****  
        8'b01100000, // 1  **     
        8'b11000000, // 2 **      
        8'b11111100, // 3 ******  
        8'b11000110, // 4 **   ** 
        8'b11000110, // 5 **   ** 
        8'b01111100, // 6  *****  
        8'b00000000, // 7         
         // code x07
        8'b11111110, // 0 ******* 
        8'b11000110, // 1 **   ** 
        8'b00001100, // 2     **  
        8'b00011000, // 3    **   
        8'b00110000, // 4   **    
        8'b00110000, // 5   **    
        8'b00110000, // 6   **    
        8'b00000000, // 7         
         // code x08
        8'b01111000, // 0  ****   
        8'b11000100, // 1 **   *  
        8'b11100100, // 2 ***  *  
        8'b01111000, // 3  ****   
        8'b10011110, // 4 *  **** 
        8'b10000110, // 5 *    ** 
        8'b01111100, // 6  *****  
        8'b00000000, // 7         
         // code x09
        8'b01111100, // 0  *****  
        8'b11000110, // 1 **   ** 
        8'b11000110, // 2 **   ** 
        8'b01111110, // 3  ****** 
        8'b00000110, // 4      ** 
        8'b00001100, // 5     **  
        8'b01111000, // 6  ****   
        8'b00000000, // 7         
         // code x0a
        8'b00111000, // 0   ***   
        8'b01101100, // 1  ** **  
        8'b11000110, // 2 **   ** 
        8'b11000110, // 3 **   ** 
        8'b11111110, // 4 ******* 
        8'b11000110, // 5 **   ** 
        8'b11000110, // 6 **   ** 
        8'b00000000, // 7         
         // code x0b
        8'b11111100, // 0 ******  
        8'b11000110, // 1 **   ** 
        8'b11000110, // 2 **   ** 
        8'b11111100, // 3 ******  
        8'b11000110, // 4 **   ** 
        8'b11000110, // 5 **   ** 
        8'b11111100, // 6 ******  
        8'b00000000, // 7         
         // code x0c
        8'b00111100, // 0   ****  
        8'b01100110, // 1  **  ** 
        8'b11000000, // 2 **      
        8'b11000000, // 3 **      
        8'b11000000, // 4 **      
        8'b01100110, // 5  **  ** 
        8'b00111100, // 6   ****  
        8'b00000000, // 7         
         // code x0d
        8'b11111000, // 0 *****   
        8'b11001100, // 1 **  **  
        8'b11000110, // 2 **   ** 
        8'b11000110, // 3 **   ** 
        8'b11000110, // 4 **   ** 
        8'b11001100, // 5 **  **  
        8'b11111000, // 6 *****   
        8'b00000000, // 7         
         // code x0e
        8'b11111110, // 0 ******* 
        8'b11000000, // 1 **      
        8'b11000000, // 2 **      
        8'b11111100, // 3 ******  
        8'b11000000, // 4 **      
        8'b11000000, // 5 **      
        8'b11111110, // 6 ******* 
        8'b00000000, // 7         
         // code x0f
        8'b11111110, // 0 ******* 
        8'b11000000, // 1 **      
        8'b11000000, // 2 **      
        8'b11111100, // 3 ******  
        8'b11000000, // 4 **      
        8'b11000000, // 5 **      
        8'b11000000, // 6 **      
        8'b00000000, // 7         
         // code x10
        8'b00111110, // 0   ***** 
        8'b01100000, // 1  **     
        8'b11000000, // 2 **      
        8'b11001110, // 3 **  *** 
        8'b11000110, // 4 **   ** 
        8'b01100110, // 5  **  ** 
        8'b00111110, // 6   ***** 
        8'b00000000, // 7         
         // code x11
        8'b11000110, // 0 **   ** 
        8'b11000110, // 1 **   ** 
        8'b11000110, // 2 **   ** 
        8'b11111110, // 3 ******* 
        8'b11000110, // 4 **   ** 
        8'b11000110, // 5 **   ** 
        8'b11000110, // 6 **   ** 
        8'b00000000, // 7         
         // code x12
        8'b11111100, // 0 ******  
        8'b00110000, // 1   **    
        8'b00110000, // 2   **    
        8'b00110000, // 3   **    
        8'b00110000, // 4   **    
        8'b00110000, // 5   **    
        8'b11111100, // 6 ******  
        8'b00000000, // 7         
         // code x13
        8'b00000110, // 0      ** 
        8'b00000110, // 1      ** 
        8'b00000110, // 2      ** 
        8'b00000110, // 3      ** 
        8'b00000110, // 4      ** 
        8'b11000110, // 5 **   ** 
        8'b01111100, // 6  *****  
        8'b00000000, // 7         
         // code x14
        8'b11000110, // 0 **   ** 
        8'b11001100, // 1 **  **  
        8'b11011000, // 2 ** **   
        8'b11110000, // 3 ****    
        8'b11111000, // 4 *****   
        8'b11011100, // 5 ** ***  
        8'b11001110, // 6 **  *** 
        8'b00000000, // 7         
         // code x15
        8'b11000000, // 0 **      
        8'b11000000, // 1 **      
        8'b11000000, // 2 **      
        8'b11000000, // 3 **      
        8'b11000000, // 4 **      
        8'b11000000, // 5 **      
        8'b11111110, // 6 ******* 
        8'b00000000, // 7         
         // code x16
        8'b11000110, // 0 **   ** 
        8'b11101110, // 1 *** *** 
        8'b11111110, // 2 ******* 
        8'b11111110, // 3 ******* 
        8'b11010110, // 4 ** * ** 
        8'b11000110, // 5 **   ** 
        8'b11000110, // 6 **   ** 
        8'b00000000, // 7         
         // code x17
        8'b11000110, // 0 **   ** 
        8'b11100110, // 1 ***  ** 
        8'b11110110, // 2 **** ** 
        8'b11111110, // 3 ******* 
        8'b11011110, // 4 ** **** 
        8'b11001110, // 5 **  *** 
        8'b11000110, // 6 **   ** 
        8'b00000000, // 7         
         // code x18
        8'b01111100, // 0  *****  
        8'b11000110, // 1 **   ** 
        8'b11000110, // 2 **   ** 
        8'b11000110, // 3 **   ** 
        8'b11000110, // 4 **   ** 
        8'b11000110, // 5 **   ** 
        8'b01111100, // 6  *****  
        8'b00000000, // 7         
         // code x19
        8'b11111100, // 0 ******  
        8'b11000110, // 1 **   ** 
        8'b11000110, // 2 **   ** 
        8'b11000110, // 3 **   ** 
        8'b11111100, // 4 ******  
        8'b11000000, // 5 **      
        8'b11000000, // 6 **      
        8'b00000000, // 7         
         // code x1a
        8'b01111100, // 0  *****  
        8'b11000110, // 1 **   ** 
        8'b11000110, // 2 **   ** 
        8'b11000110, // 3 **   ** 
        8'b11011110, // 4 ** **** 
        8'b11001100, // 5 **  **  
        8'b01111010, // 6  **** * 
        8'b00000000, // 7         
         // code x1b
        8'b11111100, // 0 ******  
        8'b11000110, // 1 **   ** 
        8'b11000110, // 2 **   ** 
        8'b11001100, // 3 **  **  
        8'b11111000, // 4 *****   
        8'b11011100, // 5 ** ***  
        8'b11001110, // 6 **  *** 
        8'b00000000, // 7         
         // code x1c
        8'b01111000, // 0  ****   
        8'b11001100, // 1 **  **  
        8'b11000000, // 2 **      
        8'b01111100, // 3  *****  
        8'b00000110, // 4      ** 
        8'b11000110, // 5 **   ** 
        8'b01111100, // 6  *****  
        8'b00000000, // 7         
         // code x1d
        8'b11111100, // 0 ******  
        8'b00110000, // 1   **    
        8'b00110000, // 2   **    
        8'b00110000, // 3   **    
        8'b00110000, // 4   **    
        8'b00110000, // 5   **    
        8'b00110000, // 6   **    
        8'b00000000, // 7         
         // code x1e
        8'b11000110, // 0 **   ** 
        8'b11000110, // 1 **   ** 
        8'b11000110, // 2 **   ** 
        8'b11000110, // 3 **   ** 
        8'b11000110, // 4 **   ** 
        8'b11000110, // 5 **   ** 
        8'b01111100, // 6  *****  
        8'b00000000, // 7         
         // code x1f
        8'b11000110, // 0 **   ** 
        8'b11000110, // 1 **   ** 
        8'b11000110, // 2 **   ** 
        8'b11101110, // 3 *** *** 
        8'b01111100, // 4  *****  
        8'b00111000, // 5   ***   
        8'b00010000, // 6    *    
        8'b00000000, // 7         
         // code x20
        8'b11000110, // 0 **   ** 
        8'b11000110, // 1 **   ** 
        8'b11010110, // 2 ** * ** 
        8'b11111110, // 3 ******* 
        8'b11111110, // 4 ******* 
        8'b11101110, // 5 *** *** 
        8'b11000110, // 6 **   ** 
        8'b00000000, // 7         
         // code x21
        8'b11000110, // 0 **   ** 
        8'b11101110, // 1 *** *** 
        8'b01111100, // 2  *****  
        8'b00111000, // 3   ***   
        8'b01111100, // 4  *****  
        8'b11101110, // 5 *** *** 
        8'b11000110, // 6 **   ** 
        8'b00000000, // 7         
         // code x22
        8'b11001100, // 0 **  **  
        8'b11001100, // 1 **  **  
        8'b11001100, // 2 **  **  
        8'b01111000, // 3  ****   
        8'b00110000, // 4   **    
        8'b00110000, // 5   **    
        8'b00110000, // 6   **    
        8'b00000000, // 7         
         // code x23
        8'b11111110, // 0 ******* 
        8'b00001110, // 1     *** 
        8'b00011100, // 2    ***  
        8'b00111000, // 3   ***   
        8'b01110000, // 4  ***    
        8'b11100000, // 5 ***     
        8'b11111110, // 6 ******* 
        8'b00000000, // 7         
         // code x24
        8'b00000000, // 0         
        8'b00000000, // 1         
        8'b00000000, // 2         
        8'b00000000, // 3         
        8'b00000000, // 4         
        8'b01100000, // 5  **     
        8'b01100000, // 6  **     
        8'b00000000, // 7         
         // code x25
        8'b00000000, // 0         
        8'b00000000, // 1         
        8'b00000000, // 2         
        8'b00000000, // 3         
        8'b00000000, // 4         
        8'b00011000, // 5    **   
        8'b00001000, // 6     *   
        8'b00010000, // 7    *    
         // code x26
        8'b00110000, // 0   **    
        8'b00110000, // 1   **    
        8'b00110000, // 2   **    
        8'b00110000, // 3   **    
        8'b00110000, // 4   **    
        8'b00000000, // 5         
        8'b00110000, // 6   **    
        8'b00000000, // 7         
         // code x27
        8'b00100100, // 0   *  *  
        8'b01111110, // 1  ****** 
        8'b00100100, // 2   *  *  
        8'b00100100, // 3   *  *  
        8'b01111110, // 4  ****** 
        8'b00100100, // 5   *  *  
        8'b00000000, // 6         
        8'b00000000, // 7         
         // code x28
        8'b00000000, // 0         
        8'b00000000, // 1         
        8'b00000000, // 2         
        8'b01111100, // 3  *****  
        8'b00000000, // 4         
        8'b00000000, // 5         
        8'b00000000, // 6         
        8'b00000000, // 7         
         // code x29
        8'b00000011, // 0       **
        8'b00000110, // 1      ** 
        8'b00001100, // 2     **  
        8'b00011000, // 3    **   
        8'b00110000, // 4   **    
        8'b01100000, // 5  **     
        8'b11000000, // 6 **      
        8'b00000000, // 7         
         // code x2a
        8'b00000000, // 0         
        8'b00011000, // 1    **   
        8'b00011000, // 2    **   
        8'b00000000, // 3         
        8'b00000000, // 4         
        8'b00011000, // 5    **   
        8'b00011000, // 6    **   
        8'b00000000, // 7         
         // code x2b
        8'b00000000, // 0         
        8'b00000000, // 1         
        8'b01111100, // 2  *****  
        8'b00000000, // 3         
        8'b00000000, // 4         
        8'b01111100, // 5  *****  
        8'b00000000, // 6         
        8'b00000000, // 7         
         // code x2c
        8'b00111000, // 0   ***   
        8'b01000100, // 1  *   *  
        8'b10111010, // 2 * *** * 
        8'b10100010, // 3 * *   * 
        8'b10100010, // 4 * *   * 
        8'b10111010, // 5 * *** * 
        8'b01000100, // 6  *   *  
        8'b00111000, // 7   ***   
        };

	assign data = ROM[addr];

endmodule  