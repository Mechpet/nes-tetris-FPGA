package template_pkg;

parameter [1:0] BLACK = 2'b00;
parameter [1:0] DARK = 2'b01;
parameter [1:0] LIGHT = 2'b10;
parameter [1:0] WHITE = 2'b11;

parameter [6:0] O_start = 0;
parameter [6:0] I_start = 4;
parameter [6:0] Z_start = 12;
parameter [6:0] S_start = 20;
parameter [6:0] T_start = 28;
parameter [6:0] J_start = 44;
parameter [6:0] L_start = 60;

endpackage